LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

--! This package contains the functions used in the design.
PACKAGE function_pack IS

END PACKAGE function_pack;

PACKAGE BODY function_pack IS

END PACKAGE BODY function_pack;