LIBRARY IEEE;

USE IEEE.std_logic_1164.ALL;
USE IEEE.std_logic_arith.ALL;

PACKAGE MyPackage IS

  CONSTANT MY_CONSTANT : INTEGER := 10;

  TYPE my_type IS ARRAY (0 TO 7) OF STD_LOGIC;

  FUNCTION my_function(a : STD_LOGIC; b : INTEGER) RETURN STD_LOGIC;
END PACKAGE MyPackage;

PACKAGE BODY MyPackage IS

  FUNCTION my_function(a : STD_LOGIC; b : INTEGER) RETURN STD_LOGIC IS
  BEGIN
    IF a = '1' THEN
      RETURN '0';
    ELSE
      RETURN '1';
    END IF;
  END FUNCTION;

END PACKAGE BODY MyPackage;